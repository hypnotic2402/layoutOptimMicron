* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and_dummy                                    *
* Netlisted  : Tue Jan 16 10:08:51 2024                     *
* PVS Version: 21.12-s022 Wed Feb 9 12:12:42 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_2                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_2 B_botTap D_drain_1 S_source_0 4 5
** N=5 EP=5 FDC=1
M0 D_drain_1 4 S_source_0 5 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 B_topTap D_drain_1 S_source_0 4
** N=5 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_topTap g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=101.688 scb=0.082094 scc=0.0121216 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_4 B_botTap D_drain_1 S_source_0 4
** N=4 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_botTap g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and_dummy                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and_dummy GND VCC VINA VINB VOUT VOUTNAND
** N=7 EP=6 FDC=6
X4 4 VOUTNAND 4 VINA GND nmos1v_CDNS_2 $T=1600 4400 0 0 $X=1180 $Y=3840
X5 GND 4 GND VINB GND nmos1v_CDNS_2 $T=4000 1580 0 0 $X=3580 $Y=1020
X6 VCC VOUTNAND VCC VINA pmos1v_CDNS_3 $T=1600 7600 0 0 $X=1180 $Y=7400
X7 VCC VOUTNAND VCC VINB pmos1v_CDNS_3 $T=4000 7600 0 0 $X=3580 $Y=7400
X8 VCC VOUT VCC VOUTNAND pmos1v_CDNS_3 $T=6460 7600 0 0 $X=6040 $Y=7400
X9 GND VOUT GND VOUTNAND nmos1v_CDNS_4 $T=6460 3880 0 0 $X=6040 $Y=3320
.ends and_dummy
