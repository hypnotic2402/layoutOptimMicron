* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv_dummy                                    *
* Netlisted  : Tue Jan 16 10:02:14 2024                     *
* PVS Version: 21.12-s022 Wed Feb 9 12:12:42 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_2                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_2 B_botTap D_drain_1 S_source_0 4
** N=4 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_botTap g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.10409 scb=0.000241229 scc=2.8103e-08 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 B_topTap D_drain_1 S_source_0 4
** N=5 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_topTap g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=101.688 scb=0.082094 scc=0.0121216 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_dummy                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_dummy GND VCC VIN VOUT
** N=4 EP=4 FDC=2
X0 GND VOUT GND VIN nmos1v_CDNS_2 $T=1540 1080 0 0 $X=1120 $Y=520
X1 VCC VOUT VCC VIN pmos1v_CDNS_3 $T=1540 3080 0 0 $X=1120 $Y=2880
.ends inv_dummy
