* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : design_combo_2                               *
* Netlisted  : Tue Mar 19 15:07:05 2024                     *
* PVS Version: 21.12-s022 Wed Feb 9 12:12:42 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_4 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=101.688 scb=0.082094 scc=0.0121216 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_dummy                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_dummy 1 2 3 4
** N=4 EP=4 FDC=2
X2 2 4 1 pmos1v_CDNS_4 $T=1540 3080 0 0 $X=1120 $Y=2880
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.10409 scb=0.000241229 scc=2.8103e-08 $X=1540 $Y=1080 $dt=0
.ends inv_dummy

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_5                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_5 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=75.4216 scb=0.0690683 scc=0.00879748 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nor_dummy                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nor_dummy 1 2 3 4 5
** N=6 EP=5 FDC=4
X4 3 6 1 pmos1v_CDNS_5 $T=1080 3620 0 0 $X=660 $Y=3420
X5 6 4 2 pmos1v_CDNS_5 $T=3440 2720 0 0 $X=3020 $Y=2520
M0 4 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1080 $Y=1140 $dt=0
M1 4 2 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=5.05241 scb=0.000962138 scc=1.23864e-06 $X=3440 $Y=1140 $dt=0
.ends nor_dummy

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand_dummy                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand_dummy 1 2 3 4 5
** N=6 EP=5 FDC=4
X2 3 4 1 pmos1v_CDNS_4 $T=1440 3880 0 0 $X=1020 $Y=3680
X3 3 4 2 pmos1v_CDNS_4 $T=3320 3880 0 0 $X=2900 $Y=3680
M0 4 1 6 5 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=1440 $Y=2700 $dt=0
M1 6 2 5 5 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 $X=3320 $Y=1080 $dt=0
.ends nand_dummy

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: design_combo_2                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt design_combo_2
** N=28 EP=0 FDC=56
X23 12 13 14 1 inv_dummy $T=-9380 17320 0 0 $X=-9580 $Y=17320
X24 1 13 14 2 inv_dummy $T=-3580 25610 0 0 $X=-3780 $Y=25610
X25 1 13 14 3 inv_dummy $T=170 10870 0 0 $X=-30 $Y=10870
X26 2 13 14 15 inv_dummy $T=4270 35430 0 0 $X=4070 $Y=35430
X27 3 13 14 16 inv_dummy $T=10030 1040 0 0 $X=9830 $Y=1040
X28 17 13 14 18 inv_dummy $T=25680 10870 0 0 $X=25480 $Y=10870
X29 19 13 14 5 inv_dummy $T=25680 28060 0 0 $X=25480 $Y=28060
X30 20 13 14 6 inv_dummy $T=36110 16700 0 0 $X=35910 $Y=16700
X31 6 13 14 7 inv_dummy $T=39960 24990 0 0 $X=39760 $Y=24990
X32 6 13 14 8 inv_dummy $T=43010 10250 0 0 $X=42810 $Y=10250
X33 7 13 14 9 inv_dummy $T=45480 34820 0 0 $X=45280 $Y=34820
X34 8 13 14 21 inv_dummy $T=49550 1280 0 0 $X=49350 $Y=1280
X35 22 13 14 11 inv_dummy $T=63640 27450 0 0 $X=63440 $Y=27450
X36 23 13 14 24 inv_dummy $T=65930 10250 0 0 $X=65730 $Y=10250
X37 15 4 13 19 14 nor_dummy $T=12520 27160 0 0 $X=12520 $Y=27160
X38 5 18 13 20 14 nor_dummy $T=28710 18260 0 0 $X=28710 $Y=18260
X39 9 10 13 22 14 nor_dummy $T=54560 26550 0 0 $X=54560 $Y=26550
X40 2 3 13 4 14 nand_dummy $T=8830 17750 0 0 $X=8830 $Y=17750
X41 4 16 13 17 14 nand_dummy $T=17070 10380 0 0 $X=17070 $Y=10380
X42 7 8 13 10 14 nand_dummy $T=49640 17140 0 0 $X=49640 $Y=17140
X43 10 21 13 23 14 nand_dummy $T=58230 9770 0 0 $X=58230 $Y=9770
.ends design_combo_2
