* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv3_dummy                                   *
* Netlisted  : Tue Jan 16 10:04:33 2024                     *
* PVS Version: 21.12-s022 Wed Feb 9 12:12:42 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_2                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_2 B_botTap D_drain_1 S_source_0 4
** N=4 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_botTap g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.87363 scb=0.000164669 scc=8.05949e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 B_topTap D_drain_1 S_source_0 4
** N=5 EP=4 FDC=1
M0 D_drain_1 4 S_source_0 B_topTap g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=101.688 scb=0.082094 scc=0.0121216 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv3_dummy                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv3_dummy GND VCC VIN VINB VINBB VOUT
** N=6 EP=6 FDC=6
X4 GND VINB GND VIN nmos1v_CDNS_2 $T=1400 2000 0 0 $X=980 $Y=1440
X5 GND VINBB GND VINB nmos1v_CDNS_2 $T=3080 2000 0 0 $X=2660 $Y=1440
X6 GND VOUT GND VINBB nmos1v_CDNS_2 $T=4660 2000 0 0 $X=4240 $Y=1440
X7 VCC VINB VCC VIN pmos1v_CDNS_3 $T=1400 4180 0 0 $X=980 $Y=3980
X8 VCC VINBB VCC VINB pmos1v_CDNS_3 $T=3080 4180 0 0 $X=2660 $Y=3980
X9 VCC VOUT VCC VINBB pmos1v_CDNS_3 $T=4660 4180 0 0 $X=4240 $Y=3980
.ends inv3_dummy
